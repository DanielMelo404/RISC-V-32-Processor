library verilog;
use verilog.vl_types.all;
entity MagicMemory_tb is
end MagicMemory_tb;
