library verilog;
use verilog.vl_types.all;
entity InstructionDecoder is
    generic(
        opOpImm         : vl_logic_vector(6 downto 0) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1);
        opOp            : vl_logic_vector(6 downto 0) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1);
        opLui           : vl_logic_vector(6 downto 0) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1);
        opJal           : vl_logic_vector(6 downto 0) := (Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1);
        opJalr          : vl_logic_vector(6 downto 0) := (Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1);
        opBranch        : vl_logic_vector(6 downto 0) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1);
        opLoad          : vl_logic_vector(6 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        opStore         : vl_logic_vector(6 downto 0) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1);
        opAuipc         : vl_logic_vector(6 downto 0) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1);
        fnADD           : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        fnSLL           : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi1);
        fnSLT           : vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi0);
        fnSLTU          : vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi1);
        fnXOR           : vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        fnSR            : vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi1);
        fnOR            : vl_logic_vector(2 downto 0) := (Hi1, Hi1, Hi0);
        fnAND           : vl_logic_vector(2 downto 0) := (Hi1, Hi1, Hi1);
        fnBEQ           : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        fnBNE           : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi1);
        fnBLT           : vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        fnBGE           : vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi1);
        fnBLTU          : vl_logic_vector(2 downto 0) := (Hi1, Hi1, Hi0);
        fnBGEU          : vl_logic_vector(2 downto 0) := (Hi1, Hi1, Hi1);
        fnLW            : vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi0);
        fnLB            : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        fnLH            : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi1);
        fnLBU           : vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        fnLHU           : vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi1);
        fnSW            : vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi0);
        fnSB            : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        fnSH            : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi1);
        fnJALR          : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        OP              : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        OPIMM           : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        BRANCH          : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi1, Hi0);
        LUI             : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi1, Hi1);
        JAL             : vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi0, Hi0);
        JALR            : vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi0, Hi1);
        LOAD            : vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi1, Hi0);
        STORE           : vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi1, Hi1);
        AUIPC           : vl_logic_vector(3 downto 0) := (Hi1, Hi0, Hi0, Hi0);
        Unsupported     : vl_logic_vector(3 downto 0) := (Hi1, Hi0, Hi0, Hi1);
        Add             : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        Sub             : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        \And\           : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi1, Hi0);
        \Or\            : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi1, Hi1);
        \Xor\           : vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi0, Hi0);
        Slt             : vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi0, Hi1);
        Sltu            : vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi1, Hi0);
        \Sll\           : vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi1, Hi1);
        \Srl\           : vl_logic_vector(3 downto 0) := (Hi1, Hi0, Hi0, Hi0);
        \Sra\           : vl_logic_vector(3 downto 0) := (Hi1, Hi0, Hi0, Hi1);
        aluD            : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        Eq              : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        Neq             : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        Lt              : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        Ltu             : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        Ge              : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        Geu             : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi1);
        Dbr             : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0)
    );
    port(
        inst            : in     vl_logic_vector(31 downto 0);
        iType_out       : out    vl_logic_vector(3 downto 0);
        aluFunc_out     : out    vl_logic_vector(3 downto 0);
        brFunc_out      : out    vl_logic_vector(2 downto 0);
        rdIndex_out     : out    vl_logic_vector(4 downto 0);
        werf            : out    vl_logic;
        R1Index_out     : out    vl_logic_vector(4 downto 0);
        R2Index_out     : out    vl_logic_vector(4 downto 0);
        immediate_out   : out    vl_logic_vector(31 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of opOpImm : constant is 2;
    attribute mti_svvh_generic_type of opOp : constant is 2;
    attribute mti_svvh_generic_type of opLui : constant is 2;
    attribute mti_svvh_generic_type of opJal : constant is 2;
    attribute mti_svvh_generic_type of opJalr : constant is 2;
    attribute mti_svvh_generic_type of opBranch : constant is 2;
    attribute mti_svvh_generic_type of opLoad : constant is 2;
    attribute mti_svvh_generic_type of opStore : constant is 2;
    attribute mti_svvh_generic_type of opAuipc : constant is 2;
    attribute mti_svvh_generic_type of fnADD : constant is 2;
    attribute mti_svvh_generic_type of fnSLL : constant is 2;
    attribute mti_svvh_generic_type of fnSLT : constant is 2;
    attribute mti_svvh_generic_type of fnSLTU : constant is 2;
    attribute mti_svvh_generic_type of fnXOR : constant is 2;
    attribute mti_svvh_generic_type of fnSR : constant is 2;
    attribute mti_svvh_generic_type of fnOR : constant is 2;
    attribute mti_svvh_generic_type of fnAND : constant is 2;
    attribute mti_svvh_generic_type of fnBEQ : constant is 2;
    attribute mti_svvh_generic_type of fnBNE : constant is 2;
    attribute mti_svvh_generic_type of fnBLT : constant is 2;
    attribute mti_svvh_generic_type of fnBGE : constant is 2;
    attribute mti_svvh_generic_type of fnBLTU : constant is 2;
    attribute mti_svvh_generic_type of fnBGEU : constant is 2;
    attribute mti_svvh_generic_type of fnLW : constant is 2;
    attribute mti_svvh_generic_type of fnLB : constant is 2;
    attribute mti_svvh_generic_type of fnLH : constant is 2;
    attribute mti_svvh_generic_type of fnLBU : constant is 2;
    attribute mti_svvh_generic_type of fnLHU : constant is 2;
    attribute mti_svvh_generic_type of fnSW : constant is 2;
    attribute mti_svvh_generic_type of fnSB : constant is 2;
    attribute mti_svvh_generic_type of fnSH : constant is 2;
    attribute mti_svvh_generic_type of fnJALR : constant is 2;
    attribute mti_svvh_generic_type of OP : constant is 2;
    attribute mti_svvh_generic_type of OPIMM : constant is 2;
    attribute mti_svvh_generic_type of BRANCH : constant is 2;
    attribute mti_svvh_generic_type of LUI : constant is 2;
    attribute mti_svvh_generic_type of JAL : constant is 2;
    attribute mti_svvh_generic_type of JALR : constant is 2;
    attribute mti_svvh_generic_type of LOAD : constant is 2;
    attribute mti_svvh_generic_type of STORE : constant is 2;
    attribute mti_svvh_generic_type of AUIPC : constant is 2;
    attribute mti_svvh_generic_type of Unsupported : constant is 2;
    attribute mti_svvh_generic_type of Add : constant is 2;
    attribute mti_svvh_generic_type of Sub : constant is 2;
    attribute mti_svvh_generic_type of \And\ : constant is 2;
    attribute mti_svvh_generic_type of \Or\ : constant is 2;
    attribute mti_svvh_generic_type of \Xor\ : constant is 2;
    attribute mti_svvh_generic_type of Slt : constant is 2;
    attribute mti_svvh_generic_type of Sltu : constant is 2;
    attribute mti_svvh_generic_type of \Sll\ : constant is 2;
    attribute mti_svvh_generic_type of \Srl\ : constant is 2;
    attribute mti_svvh_generic_type of \Sra\ : constant is 2;
    attribute mti_svvh_generic_type of aluD : constant is 2;
    attribute mti_svvh_generic_type of Eq : constant is 1;
    attribute mti_svvh_generic_type of Neq : constant is 1;
    attribute mti_svvh_generic_type of Lt : constant is 1;
    attribute mti_svvh_generic_type of Ltu : constant is 1;
    attribute mti_svvh_generic_type of Ge : constant is 1;
    attribute mti_svvh_generic_type of Geu : constant is 1;
    attribute mti_svvh_generic_type of Dbr : constant is 1;
end InstructionDecoder;
