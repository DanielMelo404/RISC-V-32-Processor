module InstructionDecoder_tb;
    reg [31:0] inst;
    
    wire [3:0] iType_out;
    wire [3:0] aluFunc_out;
    wire [2:0] brFunc_out;
    wire [4:0] rdIndex_out;
    wire werf;
    wire [4:0] R1Index_out;
    wire [4:0] R2Index_out;
    wire [31:0] immediate_out;


    InstructionDecoder uut(
    //INPUT
    .inst(inst),
    //OUTPUTS
    .iType_out(iType_out),
    .aluFunc_out(aluFunc_out),
    .brFunc_out(brFunc_out),
    .rdIndex_out(rdIndex_out),
    .werf(werf),
    .R1Index_out(R1Index_out),
    .R2Index_out(R2Index_out),
    .immediate_out(immediate_out)
    );

    initial begin
        
        inst = 32'b00000000010000001000000010010011; //addi x1, x1, 4//-------------------OPIMM
        #10
        inst = 32'b10010101100100100010000100010011; //slti x2, x4, 0b1001010110010
        #10
        inst = 32'b01010010100110100011010010010011; //sltiu x9, x20, 0b0101001010011
        #10
        inst = 32'b11111000001100010100001010010011; //xori  x5, x2, 0b1111100000110
        #10
        inst = 32'b00011100011011001110010010010011; //ori  x9, x25, 0b0001110001100
        #10
        inst = 32'b10101010011101100111011110010011; //andi  x15, x12, 0b1010101001110
        #10
        inst = 32'b00000000011001100001100100010011; //slli  x18, x12, 0b00110
        #10
        inst = 32'b00000001011001100101100100010011; //srli  x18, x12, 0b10110
        #10
        inst = 32'b01000000001101000101010100010011; //srai  x10, x8, 0b01110
        #10
        inst = 32'b00000000011001000000010100110011; //add  x10, x8, x6//-------------------OP
        #10
        inst = 32'b01000000011001000000010100110011; //sub  x10, x8, x6
        #10
        inst = 32'b00000000011001000001010100110011; //sll  x10, x8, x6
        #10
        inst = 32'b00000000011001000010010100110011; //slt  x10, x8, x6
        #10
        inst = 32'b00000000011001000011010100110011; //sltu  x10, x8, x6
        #10
        inst = 32'b00000000011001000100010100110011; //xor  x10, x8, x6
        #10
        inst = 32'b00000000011001000101010100110011; //srl  x10, x8, x6
        #10
        inst = 32'b01000000011001000101010100110011; //sra  x10, x8, x6
        #10
        inst = 32'b00000000011001000110010100110011; //or  x10, x8, x6
        #10
        inst = 32'b0000000001100100011101010_0110011; //and  x10, x8, x6
        #10
        inst = 32'b0000000001100100000001010_1100011; //beq x8, x6, label(10)//-------------------BRANCH
        #10
        inst = 32'b0000000001100100000101010_1100011; //bne x8, x6, label(10)
        #10
        inst = 32'b0000000001100100010001010_1100011; //blt x8, x6, label(10)
        #10
        inst = 32'b0000000001100100010101010_1100011; //bge x8, x6, label(10)
        #10
        inst = 32'b0000000_00110_01000_110_01010_1100011; //bltu x8, x6, label(10)
        #10
        inst = 32'b0000000_00110_01000_111_01010_1100011; //bgeu x8, x6, label(10)
        #10
        inst = 32'b00000000000000000001000010110111; // LUI x1, 1//-------------------LUI
        #10
        inst = 32'b00000000000000000001000011101111; // JAL x1, 20 (salta a 4096)//-------------------JAL
        #10
        inst = 32'b000000000110_01000_000_01010_1100111; //JALR  x10, offset(x8) offset de 6//-------------------JALR
        #10
        inst = 32'b000000001001_01000_010_01010_0000011; //lw  x10, offset(x8) offset de 9//-------------------LOAD
        #10
        inst = 32'b0000001_00110_01000_010_01010_0100011; //sw  x6, offset(x8) offset de 42//-------------------STORE
        #10
        $stop;
        
    end

endmodule