library verilog;
use verilog.vl_types.all;
entity addSub_fastAdd is
    generic(
        n               : integer := 1
    );
    port(
        a               : in     vl_logic_vector;
        b               : in     vl_logic_vector;
        isSub           : in     vl_logic;
        \out\           : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of n : constant is 1;
end addSub_fastAdd;
