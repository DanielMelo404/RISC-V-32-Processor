library verilog;
use verilog.vl_types.all;
entity InstructionDecoder_tb is
end InstructionDecoder_tb;
